module full_adder(input a,b,cin,output sum,carry);
  wire w1,w2;
  xor x1(sum,a,b,cin);
  and a1(w1,a,b);
  and a2(w2,b,cin);
  
  or o1(carry,w1,w2);
endmodule
